module fg_rom (	input [7:0] 	addr,
				output [151:0]	data
				);
	parameter ADDR_WIDTH = 8;
	parameter DATA_WIDTH = 152;
	logic [ADDR_WIDTH-1:0] addr_reg;

	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		//Static, x00
		 152'h0000000000000000fff9000000000000000000,
	    152'h000000000005920eeeee000000000000000000,
	    152'h00000000000111eff376000000000000000000,
	    152'h00000000000592ef4766000000000000000000,
	    152'h0000000000025e034376000000000000000000,
	    152'h0000000000bbbdc73433dc0000000000000000,
	    152'h000000000b374bdc6347bdc300000000000000,
	    152'h00000000046a741bba7671bb30000000000000,
	    152'h0000000047a674b9dc636b9c70000000000000,
	    152'h00000000476734cd9dccbddc74000000000000,
	    152'h0000000047344bbcccbbbbcb47400000085000,
	    152'h000000036a6418582225858222258222258500,
	    152'h00000003a6341298eee8991919191999591900,
	    152'h00000036344112555555591888881888881800,
	    152'h00000037a63418222222512591515151519000,
	    152'h000000437a635547a671818281818676818000,
	    152'h00000004433994367395101184254773300000,
	    152'h00000000044224473152101520000000000000,
	    152'h000000000000bcd99c9cb00192000000000000,
	    152'h000000000000bcbbdcdcbc0000000000000000,
	    152'h00000000000bcddcbccbcdc000000000000000,
	    152'h00000000000bcd9dcbbcd9dc00000000000000,
	    152'h00000000000bcd9dcbbccd9c00000000000000,
	    152'h0000000000bcd9dcb0bbccddc0000000000000,
	    152'h0000000000bcccdc000bbcc220000000000000,
	    152'h00000000001855cb0000112998000000000000,
	    152'h00000000008599200000018558000000000000,
	    152'h000000000b82528000000b188c000000000000,
	    152'h00000000bcd8880000000bcd9dc00000000000,
	    152'h00000000bcd9db0000000bbcdcb00000000000,
	    152'h00000000bbcdcb00000000bbbb100000000000,
	    152'h000000011bbbb0000000001111800000000000,
	    152'h00000001828100000000001825800000000000,
	    152'h00000001258100000000000125800000000000,
	    152'h00000018581000000000000182800000000000,
	    152'h00000015210000000000000182800000000000,
	    152'h00000011100000000000000018110000000000,
	    152'h00000125100000000000000018258000000000,
	    152'h00001259210000000000000018825280000000,
	    152'h00001111110000000000000011111110000000,
	    //Run_1, x01
	    152'h0000000000000000fffc000000000000000000,
	    152'h000000000005c40aaaaa000000000000000000,
	    152'h000000000001110ff278000000000000000000,
	    152'h00000000000aaaaf3788000000000000000000,
	    152'h000000000aa45a023278000000000000000000,
	    152'h0000000000bbed272322d00000000000000000,
	    152'h000000000722bed8223beed000000000000000,
	    152'h00000000789231bb92821bb000000000000000,
	    152'h0000000789823dce7828dcd220000000000000,
	    152'h0000000798733decddbdeed720000000000000,
	    152'h000000227333bbddbbbbddb720000006500000,
	    152'h00000028923156444565644445644445650000,
	    152'h000002797214c6aaa6cc1c1c1c1ccc5c1c0000,
	    152'h0000027333145555555c166666166666160000,
	    152'h0000022992164444445145c151515151c00000,
	    152'h00000288998553297261646161878161600000,
	    152'h0000037888cc32972c51116453772200000000,
	    152'h00000033334432821461154320000000000000,
	    152'h00000000000bdeceedbb01c400000000000000,
	    152'h00000000000bdecbbbbb000000000000000000,
	    152'h00000000000bbdbeedbb000000000000000000,
	    152'h000000000000bbdecedb000000000000000000,
	    152'h0000000000000bbdecedb00000000000000000,
	    152'h00000000000001bbdedb440000000000000000,
	    152'h000000110000011bbdb4cc4000000000000000,
	    152'h0000014611001bd1bbb4c54000000000000000,
	    152'h0000015454111ddb1b1666b000000000000000,
	    152'h0000015641ddb1dbb111dedb00000000000000,
	    152'h0000146111bbd1bb101deceb00000000000000,
	    152'h00001510011b661100bbeedbb0000000000000,
	    152'h0000161000164546000bddbb10000000000000,
	    152'h0000110000006660000bbbb160000000000000,
	    152'h00000000000000000000111646000000000000,
	    152'h00000000000000000000016456000610000000,
	    152'h00000000000000000000001645106410000000,
	    152'h00000000000000000000000161465610000000,
	    152'h000000000000000000000000165c4100000000,
	    152'h00000000000000000000000016461000000000,
	    152'h00000000000000000000000001110000000000,
	    152'h00000000000000000000000000000000000000,
	    //Run_2, x02
	    152'h0000000000000000fffa000000000000000000,
	    152'h000000000007a90ccccc000000000000000000,
	    152'h00000000000888cff134000000000000000000,
	    152'h000000000007a9cf2344000000000000000000,
	    152'h0000000000097c012134000000000000000000,
	    152'h0000000000555de31211de0000000000000000,
	    152'h00000000051325de41235de100000000000000,
	    152'h00000000024632855634385510000000000000,
	    152'h000000001464125ade4145ae30000000000000,
	    152'h00000000134312edadee5dde32000000000000,
	    152'h000000001131255eee5555e5232000000b7000,
	    152'h0000000014638b7b9997b7b99997b99997b700,
	    152'h00000001346189abcccbaa8a8a8a8aaa7a8a00,
	    152'h000000013122897777777a8bbbbb8bbbbb8b00,
	    152'h0000000116638b9999997897a878787878a000,
	    152'h00000001446647721643b8b9b8b8b434b8b000,
	    152'h000000023444aa2163178088b2972331100000,
	    152'h0000000021119921419b808790000000000000,
	    152'h0000000000005edadde55008a9000000000000,
	    152'h0000000000005edaee55500000000000000000,
	    152'h00000000000055eedde5500000000000000000,
	    152'h000000000000055edade500000000000000000,
	    152'h0000000000000055edade50000000000000000,
	    152'h00000000000000055edade5000000000000000,
	    152'h000000000000000855ee999000000000000000,
	    152'h0000000000000005888b7a7b00000000000000,
	    152'h0000000000000005588b979b00000000000000,
	    152'h000000000000005585eebbb000000000000000,
	    152'h00000000000000558edade5000000000000000,
	    152'h00000000000008585eade50000000000000000,
	    152'h000000000000088885ee500000000000000000,
	    152'h00000000000008b8b888000000000000000000,
	    152'h0000000000008b8b97b8000000000000000000,
	    152'h0000000000008b897980000000000000000000,
	    152'h0000000000008b897b00000000000000000000,
	    152'h000000000008bb8b8800000000000000000000,
	    152'h000000000008b897a980000000000000000000,
	    152'h00000000000088b97a79b00000000000000000,
	    152'h00000000000008888888800000000000000000,
	    152'h00000000000000000000000000000000000000,
	    //Run_3, x03
	    152'h0000000000000000fff4000000000000000000,
	    152'h00000000088643088888000000000000000000,
	    152'h000000000008880ffa9d000000000000000000,
	    152'h000000000006438fb9dd000000000000000000,
	    152'h000000000008880aba9d000000000000000000,
	    152'h00000000000555c7abaa000000000000000000,
	    152'h0000000000599a5c7ab5700000000000000000,
	    152'h00000000059de9b155d9a10000000000000000,
	    152'h0000000009ded9b74c7d957000000000000000,
	    152'h0000000009de9ab774c757c000000000000000,
	    152'h000000000a99bb557777577a00000000000260,
	    152'h0000000009de9a526233362623333623333626,
	    152'h0000000009de9a134288824414141414446414,
	    152'h0000000009dbb2136666666412222212222212,
	    152'h000000000b9dda123333336136416161616140,
	    152'h000000000badeed66bae9a2123212121d9d120,
	    152'h000000000ba99e44bae9a0bb112bb36a99aa00,
	    152'h0000000000bbbb33bada000b163ba000000000,
	    152'h0000000000057c4c7c75555001430000000000,
	    152'h000000000005557c7c57cc7555000000000000,
	    152'h0000000000057755775cccc753300000000000,
	    152'h0000000000057cc75555777534630000000000,
	    152'h0000000000057c4c7555555136620000000000,
	    152'h0000000000057c4c7500551112250000000000,
	    152'h0000000000577c47500000157c750000000000,
	    152'h000000000057c4c750000057cc500000000000,
	    152'h000000000057c4750000055777500000000000,
	    152'h00000000001133350000011111000000000000,
	    152'h00000000051364620000012362000000000000,
	    152'h00000000577236320000013620000000000000,
	    152'h000000057c4721200000012300000000000000,
	    152'h0000000574c751000000121100000000000000,
	    152'h00000001577510000000123620000000000000,
	    152'h00000012111100000000112363000000000000,
	    152'h00000013431000000000001111100000000000,
	    152'h00000136210000000000000000000000000000,
	    152'h00001211000000000000000000000000000000,
	    152'h00001346200000000000000000000000000000,
	    152'h00001234632000000000000000000000000000,
	    152'h00000111111000000000000000000000000000,
	    //Run_4, x04
	    152'h0000000000000000fffb000000000000000000,
	    152'h000000000008b90ccccc000000000000000000,
	    152'h00000000000777cff134000000000000000000,
	    152'h000000000008b9cf2344000000000000000000,
	    152'h0000000000098c012134000000000000000000,
	    152'h0000000000555de31211de0000000000000000,
	    152'h00000000051325de41235de100000000000000,
	    152'h00000000024632755634375510000000000000,
	    152'h000000001464125bde4145be30000000000000,
	    152'h00000000134312edbdee5dde32000000000000,
	    152'h000000001131255eee5555e5232000000a8000,
	    152'h0000000014637a8a9998a8a99998a99998a800,
	    152'h00000001346179bacccabb7b7b7b7bbb8b7b00,
	    152'h000000013122798888888b7aaaaa7aaaaa7a00,
	    152'h0000000116637a9999998798b787878787b000,
	    152'h00000001446648821643a7a9a7a7a434a7a000,
	    152'h000000023444bb2163187077a2982331100000,
	    152'h0000000021119921419a707890000000000000,
	    152'h0000000000005edbdde55007b9000000000000,
	    152'h0000000000005edbde55500000000000000000,
	    152'h00000000000055e5ebde550000000000000000,
	    152'h000000000000055eddbbde5000000000000000,
	    152'h0000000000000055edddbde500000000000000,
	    152'h000000000000000775edde5890000000000000,
	    152'h00000000000000055777778ba0000000000000,
	    152'h000000000000007775eb5798a0000000000000,
	    152'h000000000000778b75edde7a00000000000000,
	    152'h0000000000079a99875ee55000000000000000,
	    152'h000000000007ba777775500000000000000000,
	    152'h0000000000789755ee50000000000000000000,
	    152'h000000000079a7777500000000000000000000,
	    152'h00000000007977a9a700000000000000000000,
	    152'h00000000007a079a7000000000000000000000,
	    152'h0000000000777a9a7000000000000000000000,
	    152'h0000000000007aa70000000000000000000000,
	    152'h000000000007a7770000000000000000000000,
	    152'h000000000007a98a7000000000000000000000,
	    152'h0000000000077a989a70000000000000000000,
	    152'h00000000000007777770000000000000000000,
	    152'h00000000000000000000000000000000000000,
	    //Shoot_1, x05
	    152'h000000000000b000fffa000000000000000000,
	    152'h000000000b08ab0bbbbb000000000000000000,
	    152'h0000000000bb33bff157000000000000000000,
	    152'h000000000008bb0f2577000000000000000000,
	    152'h00000000000689012157000000000000000000,
	    152'h0000000000ccced51211ed0000000000000000,
	    152'h000000000c152ced7125ced100000000000000,
	    152'h000000000147523cc45753cc00000000000000,
	    152'h00000000247512caed717cad10000000000000,
	    152'h0000000027512cdeaeddceed20000000000000,
	    152'h000000025122cccdddccccdc50000000980000,
	    152'h00000014752398966689896666896666898000,
	    152'h0000014751236a74447aa3a3a3a3aaa8a3a000,
	    152'h00000151223368888888a39999939999939000,
	    152'h00000254712396666668368a383838383a0000,
	    152'h00000215471882547539396939397579390000,
	    152'h0000002211aa2175133a833926825511000000,
	    152'h0000000022662251d336938600000000000000,
	    152'h0000000000000cdeaadadc3a60000000000000,
	    152'h0000000000000cdccededcd000000000000000,
	    152'h000000000000cdeedcddcded00000000000000,
	    152'h000000000000cdeaedccdeaed0000000000000,
	    152'h000000000000cdeaedccddead0000000000000,
	    152'h00000000000cdeaedc0ccddeed000000000000,
	    152'h00000000000cddded000ccdd66000000000000,
	    152'h000000000003988dc0000336aa900000000000,
	    152'h0000000000098aa60000003988900000000000,
	    152'h0000000000c96869000000c399d00000000000,
	    152'h000000000cde9990000000cdeaed0000000000,
	    152'h000000000cdeaec0000000ccdedc0000000000,
	    152'h000000000ccdedc00000000cccc30000000000,
	    152'h0000000033cccc000000000333390000000000,
	    152'h00000000396930000000000396890000000000,
	    152'h00000000368930000000000036890000000000,
	    152'h00000003989300000000000039690000000000,
	    152'h00000003693000000000000039690000000000,
	    152'h00000003330000000000000003933000000000,
	    152'h00000036830000000000000003968900000000,
	    152'h00000368a63000000000000003996869000000,
	    152'h00000333333000000000000003333333000000,
		 
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000,
		 152'h00000000000000000000000000000000000000
				 
	    //shoot_2, x06
		 /*
	    168'h000000000000b000fffa000000000000000000,
	    168'h000000000b08ab0bbbbb000000000000000000,
	    168'h0000000000bb33bff157000000000000000000,
	    168'h000000000008bb0f2577000000000000000000,
	    168'h00000000000689012157000000000000000000,
	    168'h0000000000ccced51211ed0000000000000000,
	    168'h000000000c152ced7125ced100000000000000,
	    168'h000000000147523cc45753cc00000000000000,
	    168'h00000000247512caed717cad10000000000000,
	    168'h0000000027512cdeaeddceed20000000000000,
	    168'h000000025122cccdddccccdc50000000980000,
	    168'h00000014752398966689896666896666816000,
	    168'h0000014751236a74447aa3a3a3a3aa16161000,
	    168'h00000151223368888888a39999939999916000,
	    168'h00000254712396666668368a383838383a0000,
	    168'h00000215471882547539396939397579390000,
	    168'h0000002211aa2175133a833926825511000000,
	    168'h0000000022662251d336938600000000000000,
	    168'h0000000000000cdeaadadc3a60000000000000,
	    168'h0000000000000cdccededcd000000000000000,
	    168'h000000000000cdeedcddcded00000000000000,
	    168'h000000000000cdeaedccdeaed0000000000000,
	    168'h000000000000cdeaedccddead0000000000000,
	    168'h00000000000cdeaedc0ccddeed000000000000,
	    168'h00000000000cddded000ccdd66000000000000,
	    168'h000000000003988dc0000336aa900000000000,
	    168'h0000000000098aa60000003988900000000000,
	    168'h0000000000c96869000000c399d00000000000,
	    168'h000000000cde9990000000cdeaed0000000000,
	    168'h000000000cdeaec0000000ccdedc0000000000,
	    168'h000000000ccdedc00000000cccc30000000000,
	    168'h0000000033cccc000000000333390000000000,
	    168'h00000000396930000000000396890000000000,
	    168'h00000000368930000000000036890000000000,
	    168'h00000003989300000000000039690000000000,
	    168'h00000003693000000000000039690000000000,
	    168'h00000003330000000000000003933000000000,
	    168'h00000036830000000000000003968900000000,
	    168'h00000368a63000000000000003996869000000,
	    168'h00000333333000000000000003333333000000
		 */
	    };
    assign data = ROM[addr];

endmodule







// Width: 253
// Height: 212
// Total colors: 5
// Index and RGB values are: 
// 0:0 0 0
// 1:0 130 198
// 2:206 203 206
// 3:255 251 255
// 4:0 73 8

module background_rom( input [7:0]	addr,
					   output [1011:0] data
					   );
	parameter ADDR_WIDTH = 8;
	parameter DATA_WIDTH = 1012;
	logic [ADDR_WIDTH-1:0] addr_reg;

	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000002000000000000000000000000000000020000000000000000000000000000000000000000000000000000000200000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000030000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000002000000000000000000000000000000020000000000000002000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000020000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000030000000000000000000000000000000000000000000000000000000000000003000000000000000000000000000000030000000000000000000000000000000300000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000002000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000020000000000000000000000000000000200000000000000000000000000000002000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000010000000000000003000000000000000000000000000000030000000000000000000000000000000300000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000002000000000000000200000000000000000000000000000002000000000000000000000000000000020000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000030000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000300000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000010111111000000001111111111111111000000000000000000000000000000001011111100000000111111111111111100000000000000000000000000000000101111110000000011111111111111110000000000000000000000000000000010111111000000001111111111111,
	    1012'h1110000000000000000000000000111122222222000011112222222222222222111000000000000000000000000011112222222200001111222222222222222211100000000000000000000000001111222222220000111122222222222222221110000000000000000000000000111122222222000011112222222222222,
	    1012'h2222201111111111111111110011222222222333001122222222222222222222222220111111111111111111001122222222233300112222222222222222222222222011111111111111111100112222222223330011222222222222222222222222201111111111111111110011222222222333001122222222222222222,
	    1012'h2231011222222222222222221021122223333310102112222222222222222222223101122222222222222222102112222333331010211222222222222222222222310112222222222222222210211222233333101021122222222222222222222231011222222222222222221021122223333310102112222222222222222,
	    1012'h2310022222222222222222222211011333211022221101133322222222222222231002222222222222222222221101133321102222110113332222222222222223100222222222222222222222110113332110222211011333222222222222222310022222222222222222222211011333211022221101133322222222222,
	    1012'h3100222222222222222222221222210120002222122221011111332222222222310022222222222222222222122221012000222212222101111133222222222231002222222222222222222212222101200022221222210111113322222222223100222222222222222222221222210120002222122221011111332222222,
	    1012'h1102222222222222222222222222222112222222222222211111112111333321110222222222222222222222222222211222222222222221111111211133332111022222222222222222222222222221122222222222222111111121113333211102222222222222222222222222222112222222222222211111112111333,
	    1012'h1022222302222221022222211222222122222222122222212212001100000011102222230222222102222221122222212222222212222221221200110000001110222223022222210222222112222221222222221222222122120011000000111022222302222221022222211222222122222222122222212212001100000,
	    1012'h1222122230222222222222222222111012221222302222222222222222221110122212223022222222222222222211101222122230222222222222222222111012221222302222222222222222221110122212223022222222222222222211101222122230222222222222222222111012221222302222222222222222221,
	    1012'h0322222220022222222222222223211003222222200222222222222222232110032222222002222222222222222321100322222220022222222222222223211003222222200222222222222222232110032222222002222222222222222321100322222220022222222222222223211003222222200222222222222222232,
	    1012'h0123222222222222222222222232111001232222222222222222222222321110012322222222222222222222223211100123222222222222222222222232111001232222222222222222222222321110012322222222222222222222223211100123222222222222222222222232111001232222222222222222222222321,
	    1012'h0112332222222222222222222311111001123322222222222222222223111110011233222222222222222222231111100112332222222222222222222311111001123322222222222222222223111110011233222222222222222222231111100112332222222222222222222311111001123322222222222222222223111,
	    1012'h0111112232222222222223333121111001111122322222222222233331211110011111223222222222222333312111100111112232222222222223333121111001111122322222222222233331211110011111223222222222222333312111100111112232222222222223333121111001111122322222222222233331211,
	    1012'h0111111111213333333333322221111001111111112133333333333222211110011111111121333333333332222111100111111111213333333333322221111001111111112133333333333222211110011111111121333333333332222111100111111111213333333333322221111001111111112133333333333222211,
	    1012'h0111111112222222233332233221111001111111122222222333322332211110011111111222222223333223322111100111111112222222233332233221111001111111122222222333322332211110011111111222222223333223322111100111111112222222233332233221111001111111122222222333322332211,
	    1012'h0111111222222233132333333322111001111112222222331323333333221110011111122222223313233333332211100111111222222233132333333322111001111112222222331323333333221110011111122222223313233333332211100111111222222233132333333322111001111112222222331323333333221,
	    1012'h1120111222312222233233332222211011201112223122222332333322222110112011122231222223323333222221101120111222312222233233332222211011201112223122222332333322222110112011122231222223323333222221101120111222312222233233332222211011201112223122222332333322222,
	    1012'h1110111122332233233333332232211011101111223322332333333322322110111011112233223323333333223221101110111122332233233333332232211011101111223322332333333322322110111011112233223323333333223221101110111122332233233333332232211011101111223322332333333322322,
	    1012'h1112011122222332332333333222110111120111222223323323333332221101111201112222233233233333322211011112011122222332332333333222110111120111222223323323333332221101111201112222233233233333322211011112011122222332332333333222110111120111222223323323333332221,
	    1012'h2111211112222222233333332221001221112111122222222333333322210012211121111222222223333333222100122111211112222222233333332221001221112111122222222333333322210012211121111222222223333333222100122111211112222222233333332221001221112111122222222333333322210,
	    1012'h2211111112222222333333322110012222111111122222223333333221100122221111111222222233333332211001222211111112222222333333322110012222111111122222223333333221100122221111111222222233333332211001222211111112222222333333322110012222111111122222223333333221100,
	    1012'h2222100112222232233333211232101222221001122222322333332112321012222210011222223223333321123210122222100112222232233333211232101222221001122222322333332112321012222210011222223223333321123210122222100112222232233333211232101222221001122222322333332112321,
	    1012'h2222212111222023333311112333210122222121112220233333111123332101222221211122202333331111233321012222212111222023333311112333210122222121112220233333111123332101222221211122202333331111233321012222212111222023333311112333210122222121112220233333111123332,
	    1012'h0211122210011101221112223333321002111222100111012211122233333210021112221001110122111222333332100211122210011101221112223333321002111222100111012211122233333210021112221001110122111222333332100211122210011101221112223333321002111222100111012211122233333,
	    1012'h0111222201122310111122333332310101112222011223101111223333323101011122220112231011112233333231010111222201122310111122333332310101112222011223101111223333323101011122220112231011112233333231010111222201122310111122333332310101112222011223101111223333323,
	    1012'h0113222202222321012233333233201101132222022223210122333332332011011322220222232101223333323320110113222202222321012233333233201101132222022223210122333332332011011322220222232101223333323320110113222202222321012233333233201101132222022223210122333332332,
	    1012'h0112222022223322100232333322111101122220222233221002323333221111011222202222332210023233332211110112222022223322100232333322111101122220222233221002323333221111011222202222332210023233332211110112222022223322100232333322111101122220222233221002323333221,
	    1012'h0111220222223323101133323231012301112202222233231011333232310123011122022222332310113332323101230111220222223323101133323231012301112202222233231011333232310123011122022222332310113332323101230111220222223323101133323231012301112202222233231011333232310,
	    1012'h2111200222233332210102332321222321112002222333322101023323212223211120022223333221010233232122232111200222233332210102332321222321112002222333322101023323212223211120022223333221010233232122232111200222233332210102332321222321112002222333322101023323212,
	    1012'h2112002222233232311011233210223221120022222332323110112332102232211200222223323231101123321022322112002222233232311011233210223221120022222332323110112332102232211200222223323231101123321022322112002222233232311011233210223221120022222332323110112332102,
	    1012'h2210022122133323121101132102233222100221221333231211011321022332221002212213332312110113210223322210022122133323121101132102233222100221221333231211011321022332221002212213332312110113210223322210022122133323121101132102233222100221221333231211011321022,
	    1012'h2200222322333232321110112022232222002223223332323211101120222322220022232233323232111011202223222200222322333232321110112022232222002223223332323211101120222322220022232233323232111011202223222200222322333232321110112022232222002223223332323211101120222,
	    1012'h2220111212333313222110111011122222201112123333132221101110111222222011121233331322211011101112222220111212333313222110111011122222201112123333132221101110111222222011121233331322211011101112222220111212333313222110111011122222201112123333132221101110111,
	    1012'h2222011111133332332210010011122222220111111333323322100100111222222201111113333233221001001112222222011111133332332210010011122222220111111333323322100100111222222201111113333233221001001112222222011111133332332210010011122222220111111333323322100100111,
	    1012'h2222011111113322322210000001112222220111111133223222100000011122222201111111332232221000000111222222011111113322322210000001112222220111111133223222100000011122222201111111332232221000000111222222011111113322322210000001112222220111111133223222100000011,
	    1012'h2222000111112333233210011110111222220001111123332332100111101112222200011111233323321001111011122222000111112333233210011110111222220001111123332332100111101112222200011111233323321001111011122222000111112333233210011110111222220001111123332332100111101,
	    1012'h2220111011111232322210122211011122201110111112323222101222110111222011101111123232221012221101112220111011111232322210122211011122201110111112323222101222110111222011101111123232221012221101112220111011111232322210122211011122201110111112323222101222110,
	    1012'h1201222201111123232101222321101112012222011111232321012223211011120122220111112323210122232110111201222201111123232101222321101112012222011111232321012223211011120122220111112323210122232110111201222201111123232101222321101112012222011111232321012223211,
	    1012'h1012223210111112221012223222100110122232101111122210122232221001101222321011111222101222322210011012223210111112221012223222100110122232101111122210122232221001101222321011111222101222322210011012223210111112221012223222100110122232101111122210122232221,
	    1012'h1122232210111111210122233222110011222322101111112101222332221100112223221011111121012223322211001122232210111111210122233222110011222322101111112101222332221100112223221011111121012223322211001122232210111111210122233222110011222322101111112101222332221,
	    1012'h1322322211111111101222332222210013223222111111111012223322222100132232221111111110122233222221001322322211111111101222332222210013223222111111111012223322222100132232221111111110122233222221001322322211111111101222332222210013223222111111111012223322222,
	    1012'h1133222211000000012211322221221011332222110000000122113222212210113322221100000001221132222122101133222211000000012211322221221011332222110000000122113222212210113322221100000001221132222122101133222211000000012211322221221011332222110000000122113222212,
	    1012'h0113222210111110021112322123221001132222101111100211123221232210011322221011111002111232212322100113222210111110021112322123221001132222101111100211123221232210011322221011111002111232212322100113222210111110021112322123221001132222101111100211123221232,
	    1012'h0113222101112221011111232322222101132221011122210111112323222221011322210111222101111123232222210113222101112221011111232322222101132221011122210111112323222221011322210111222101111123232222210113222101112221011111232322222101132221011122210111112323222,
	    1012'h0111321011121223101011132222222101113210111212231010111322222221011132101112122310101113222222210111321011121223101011132222222101113210111212231010111322222221011132101112122310101113222222210111321011121223101011132222222101113210111212231010111322222,
	    1012'h0111311111122222210211112222222201113111111222222102111122222222011131111112222221021111222222220111311111122222210211112222222201113111111222222102111122222222011131111112222221021111222222220111311111122222210211112222222201113111111222222102111122222,
	    1012'h0011101111222232221011113222222200111011112222322210111132222222001110111122223222101111322222220011101111222232221011113222222200111011112222322210111132222222001110111122223222101111322222220011101111222232221011113222222200111011112222322210111132222,
	    1012'h0010011212122332222011111222222000100112121223322220111112222220001001121212233222201111122222200010011212122332222011111222222000100112121223322220111112222220001001121212233222201111122222200010011212122332222011111222222000100112121223322220111112222,
	    1012'h1011122211223323222110111111111110111222112233232221101111111111101112221122332322211011111111111011122211223323222110111111111110111222112233232221101111111111101112221122332322211011111111111011122211223323222110111111111110111222112233232221101111111,
	    1012'h0011122223233232332210011100000000111222232332323322100111000000001112222323323233221001110000000011122223233232332210011100000000111222232332323322100111000000001112222323323233221001110000000011122223233232332210011100000000111222232332323322100111000,
	    1012'h0001112211333322322210001011111000011122113333223222100010111110000111221133332232221000101111100001112211333322322210001011111000011122113333223222100010111110000111221133332232221000101111100001112211333322322210001011111000011122113333223222100010111,
	    1012'h1110111211131232233210010111222111101112111312322332100101112221111011121113123223321001011122211110111211131232233210010111222111101112111312322332100101112221111011121113123223321001011122211110111211131232233210010111222111101112111312322332100101112,
	    1012'h2211011111133212322210121112122322110111111332123222101211121223221101111113321232221012111212232211011111133212322210121112122322110111111332123222101211121223221101111113321232221012111212232211011111133212322210121112122322110111111332123222101211121,
	    1012'h2321101111123232232101221112222223211011111232322321012211122222232110111112323223210122111222222321101111123232232101221112222223211011111232322321012211122222232110111112323223210122111222222321101111123232232101221112222223211011111232322321012211122,
	    1012'h3222100111132222221012221122223232221001111322222210122211222232322210011113222222101222112222323222100111132222221012221122223232221001111322222210122211222232322210011113222222101222112222323222100111132222221012221122223232221001111322222210122211222,
	    1012'h3222110011112221210122231212233232221100111122212101222312122332322211001111222121012223121223323222110011112221210122231212233232221100111122212101222312122332322211001111222121012223121223323222110011112221210122231212233232221100111122212101222312122,
	    1012'h2221112120012332222111212001233222211121200123322221112120012332222111212001233222211121200123322221112120012332222111212001233222211121200123322221112120012332222111212001233222211121200123322221112120012332222111212001233222211121200123322221112120012,
	    1012'h2221011210002322222101121000232222210112100023222221011210002322222101121000232222210112100023222221011210002322222101121000232222210112100023222221011210002322222101121000232222210112100023222221011210002322222101121000232222210112100023222221011210002,
	    1012'h2211001111000222221100111100022222110011110002222211001111000222221100111100022222110011110002222211001111000222221100111100022222110011110002222211001111000222221100111100022222110011110002222211001111000222221100111100022222110011110002222211001111000,
	    1012'h2110000000110022211000000011002221100000001100222110000000110022211000000011002221100000001100222110000000110022211000000011002221100000001100222110000000110022211000000011002221100000001100222110000000110022211000000011002221100000001100222110000000110,
	    1012'h1100000000011001110000000001100111000000000110011100000000011001110000000001100111000000000110011100000000011001110000000001100111000000000110011100000000011001110000000001100111000000000110011100000000011001110000000001100111000000000110011100000000011,
	    1012'h0000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	    1012'h3000000000000000000000000000000330000000000000000000000000000003300000000000000000000000000000033000000000000000000000000000000330000000000000000000000000000003300000000000000000000000000000033000000000000000000000000000000330000000000000000000000000000,
	    1012'h3000000000000000000000000000000330000000000000000000000000000003300000000000000000000000000000033000000000000000000000000000000330000000000000000000000000000003300000000000000000000000000000033000000000000000000000000000000330000000000000000000000000000,
	    1012'h2300000000000000000000000000002223000000000000000000000000000022230000000000000000000000000000222300000000000000000000000000002223000000000000000000000000000022230000000000000000000000000000222300000000000000000000000000002223000000000000000000000000000,
	    1012'h2300000000000000000000000000030023000000000000000000000000000300230000000000000000000000000003002300000000000000000000000000030023000000000000000000000000000300230000000000000000000000000003002300000000000000000000000000030023000000000000000000000000000,
	    1012'h2330000000000000000000000000023023300000000000000000000000000230233000000000000000000000000002302330000000000000000000000000023023300000000000000000000000000230233000000000000000000000000002302330000000000000000000000000023023300000000000000000000000000,
	    1012'h0233000000000000000000000000220002330000000000000000000000002200023300000000000000000000000022000233000000000000000000000000220002330000000000000000000000002200023300000000000000000000000022000233000000000000000000000000220002330000000000000000000000002,
	    1012'h0002330000000000000000000330002000023300000000000000000003300020000233000000000000000000033000200002330000000000000000000330002000023300000000000000000003300020000233000000000000000000033000200002330000000000000000000330002000023300000000000000000003300,
	    1012'h3000000000000000000000000000020330000000000000000000000000000203300000000000000000000000000002033000000000000000000000000000020330000000000000000000000000000203300000000000000000000000000002033000000000000000000000000000020330000000000000000000000000000,
	    1012'h3300022000000003300000002000003233000220000000033000000020000032330002200000000330000000200000323300022000000003300000002000003233000220000000033000000020000032330002200000000330000000200000323300022000000003300000002000003233000220000000033000000020000,
	    1012'h2330000000000003330000000022432023300000000000033300000000224320233000000000000333000000002243202330000000000003330000000022432023300000000000033300000000224320233000000000000333000000002243202330000000000003330000000022432023300000000000033300000000224,
	    1012'h0223330000000022323000000000032002233300000000223230000000000320022333000000002232300000000003200223330000000022323000000000032002233300000000223230000000000320022333000000002232300000000003200223330000000022323000000000032002233300000000223230000000000,
	    1012'h0302003300000300403300003000320003020033000003004033000030003200030200330000030040330000300032000302003300000300403300003000320003020033000003004033000030003200030200330000030040330000300032000302003300000300403300003000320003020033000003004033000030003,
	    1012'h3000224000000230300300000002220330002240000002303003000000022203300022400000023030030000000222033000224000000230300300000002220330002240000002303003000000022203300022400000023030030000000222033000224000000230300300000002220330002240000002303003000000022,
	    1012'h3300000000002200333033002022000033000000000022003330330020220000330000000000220033303300202200003300000000002200333033002022000033000000000022003330330020220000330000000000220033303300202200003300000000002200333033002022000033000000000022003330330020220,
	    1012'h2232333003300020023300000000000022323330033000200233000000000000223233300330002002330000000000002232333003300020023300000000000022323330033000200233000000000000223233300330002002330000000000002232333003300020023300000000000022323330033000200233000000000,
	    1012'h2002220000000203002233000000000020022200000002030022330000000000200222000000020300223300000000002002220000000203002233000000000020022200000002030022330000000000200222000000020300223300000000002002220000000203002233000000000020022200000002030022330000000,
	    1012'h0002000000033243430044432004002000020000000332434300444320040020000200000003324343004443200400200002000000033243430044432004002000020000000332434300444320040020000200000003324343004443200400200002000000033243430044432004002000020000000332434300444320040,
	    1012'h2000020000332233233003440020032420000200003322332330034400200324200002000033223323300344002003242000020000332233233003440020032420000200003322332330034400200324200002000033223323300344002003242000020000332233233003440020032420000200003322332330034400200
	    };

	    assign data = ROM[addr];

endmodule
	   


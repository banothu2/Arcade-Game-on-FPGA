module figure_rom(input [4:0]	addr,
						output [20:0] data);
	parameter ADDR_WIDTH = 5;
	parameter DATA_WIDTH = 21;
	logic [ADDR_WIDTH-1:0] addr_reg;

	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000,
		21'b000000000000000000000
		};
		
	assign data = ROM[addr];
endmodule
